module my_jtd(
 input pka_1or2m_gck,
 input start_flag,
 input[31:0] Preamble, //为了循环所以用32位的，并非preamble是32位的。
 input rst_n,
 
 input[2:0] BLE_TYPE,
 input BLE_ADV_STATE,
 input BLE_TX_RX_EN,
 //input reg BLE_WHITEN_EN,
 input[6:0] BLE_WHITEN_INIT,
 input[23:0] BLE_CRC_INIT,
 input[31:0] BLE_ACC_ADDR, 
 input[15:0] BLE_ADV_HEADER,
 input[15:0] BLE_DATA_HEADER,
 input[1:0] BLE_CI,
 input[2:0] BLE_TERM1,
 input[2:0] BLE_TERM2,
 
 input[6:0] ram_a1,
 //input[31:0] ram_d1,
 inout[31:0] ram_d1,
 input ram_cs1,
 input ram_we1,
 input ram_oe1,

 output reg r_fsm_data
 );
 
 reg[3:0] current_state,next_state,r_cnt_cnt;
 reg[4:0] r_cnt;
 reg[7:0] r_bytes;
 reg[31:0] r_tx_shift_reg;
 reg[31:0] PAYLOAD;
 reg[6:0] RAM_A2;
 reg RAM_CS2,RAM_WEN2,RAM_OE2;
 reg r_switch_crc,r_crc_init,r_switch_dwh,tx_fsm_finished;
 reg r_rst_tx_reg; 
 
// wire[4:0] r_count;
// wire[3:0] r_cnt_count;
 wire[31:0] ram_d2;
 wire[6:0] ram_a2;
 wire ram_cs2,ram_we2,ram_oe2;
 wire switch_crc,crc_init,switch_dwh;
 wire r_rst_tx;
 
 parameter[3:0] s_idle=4'b0000,s_tx_preamble=4'b0001,s_tx_access=4'b0010,s_tx_ci=4'b0011,s_tx_term1=4'b0100,s_tx_pdu_header=4'b0101,s_tx_pdu_payload=4'b0110,s_wait_crc=4'b0111,s_tx_term2=4'b1000,s_end=4'b1001,s_reset=4'b1010;
 
 my_ram u2(.clk(pka_1or2m_gck),.a1(ram_a1),.d1(ram_d1),.we1(ram_we1),.cs1(ram_cs1),.oe1(ram_oe1),.a2(ram_a2),.d2(ram_d2),.we2(ram_we2),.cs2(ram_cs2),.oe2(ram_oe2));

assign r_rst_tx = r_rst_tx_reg;
assign ram_a2 = RAM_A2;
assign ram_cs2 = RAM_CS2;
assign ram_we2 = RAM_WEN2;
assign ram_oe2 = RAM_OE2;
assign switch_crc = r_switch_crc;
assign crc_init = r_crc_init;
assign switch_dwh = r_switch_dwh;
//assign r_count = r_cnt;
//assign r_cnt_count=r_cnt_cnt;

always@(*) 
 begin
    case(current_state)
	  s_idle: 
	    begin
		   r_fsm_data=1'b0;
         r_cnt=5'b0;
			r_cnt_cnt=4'b0;
			//if(r_tx_en)//发送使能有效，标志着发送数据准备完成
			if(BLE_TX_RX_EN) //发送使能应该在ram的payload以及preamble、header寄存器初始化，重要的就是在于ram
			//r_bytes=根据BLE_ADV_STATE的状态把当前要发送的payload的length赋值
			  begin
               r_rst_tx_reg=0;
					//注意此时默认header是16位，且只有连接和广播两种类型。
					if(BLE_ADV_STATE)    r_bytes=BLE_DATA_HEADER[15:8];
					else                 r_bytes=BLE_ADV_HEADER[15:8]; //r_bytes=length
			      
					if(start_flag)//起始时刻到来，在发送时隙的起始点或 150us 帧间隔来临
			       begin
				     r_tx_shift_reg[31:0]=Preamble[31:0];
				     next_state=s_tx_preamble;
				     r_switch_crc=1'b1;
				    end //文献：状态跳转时，需要把状态机的输出使能信号置为有效状态，同时把 CRC 模块的使能信号也置为有效状态。
				   else  next_state=s_idle;
			  end
			else next_state=s_idle;  
	    end 
     s_tx_preamble: //公共部分
	    begin
		   r_fsm_data=r_tx_shift_reg[0];  //发送数据流r_fsm_data
			r_tx_shift_reg={1'b0, r_tx_shift_reg[31:1]}; //移位
			//r_tx_shift_reg={r_tx_shift_reg[0], r_tx_shift_reg[31:1]};  
			if(BLE_TYPE==3'b010)//如果发送报文为 2Mbps 非编码类型，则在 r_cnt 第二次计数到 7 时，也就是preamble是2 octets
			  begin
			    if(r_cnt==5'd7) 
				    begin
					   r_cnt_cnt=r_cnt_cnt+4'd1;
						r_cnt=0;
					   if(r_cnt_cnt==4'd2) 
						  begin
						   r_cnt_cnt=0;
						   r_tx_shift_reg=BLE_ACC_ADDR[31:0]; 
						   next_state=s_tx_access;
						  end
						else next_state=s_tx_preamble; 
				    end
				 else next_state=s_tx_preamble;
				end
			else if(BLE_TYPE==3'b100) //如果发送报文为 1Mbps 编码类型，则在 r_cnt 第十次计数到 7 时，也就是preamble是10 octets
			  begin
			    if(r_cnt==5'd7) 
				   begin
					   r_cnt=0;
						r_cnt_cnt=r_cnt_cnt+4'd1;
					   if(r_cnt_cnt==5'd10) 
						  begin
						   r_cnt_cnt=0;
						   r_tx_shift_reg=BLE_ACC_ADDR[31:0]; 
						   next_state=s_tx_access;
						  end
						else next_state=s_tx_preamble;
				   end
				 else next_state=s_tx_preamble;
				end	
         else	//其他类型时，均在 r_cnt第一次计数到 7 时
           begin
			    if(r_cnt==5'd7) 
				   begin
					   r_cnt=0; 
						r_tx_shift_reg=BLE_ACC_ADDR[31:0]; 
						next_state=s_tx_access;
					end
				 else next_state=s_tx_preamble; 
			  end
		   r_cnt=r_cnt+5'd1;	  
       end
     s_tx_access: //公共部分
	     begin
		   r_fsm_data=r_tx_shift_reg[0];
			r_tx_shift_reg={1'b0, r_tx_shift_reg[31:1]};
         if(BLE_TYPE==3'b100) //如果发送报文为 1Mbps 编码类型，则需要把 2bits 的 CI 装载进移位寄存器，同时状态机跳转到s_tx_ci 状态
			  begin
			    if(r_cnt==5'd31)
				   begin
					   r_cnt=0;
					   r_tx_shift_reg=BLE_CI[1:0]; 
						next_state=s_tx_ci;
						r_crc_init=1'b1;//状态机跳转时，把 r_crc_init 置为 1，即对 CRC 模块进行初始化；
		            RAM_A2=7'b1111111;//同时为了方便后续对数据载荷的提取，令 TX-RAM 的地址指针指向末尾处。
				   end
				 else next_state=s_tx_access;
				end	
         else	//其他类型时，则把 16bits or 24bits （这里需要最后再解决一下，主要是数字信道的24和新的同步音频流？）的 Header 装载进移位寄存器，同时状态机跳转到 s_tx_pdu_header 状态
           begin
			    if(r_cnt==5'd31) 
				   begin
					   r_cnt=0;
						  if(BLE_ADV_STATE==0) //
						    begin
							  r_tx_shift_reg=BLE_ADV_HEADER[15:0]; 
						     next_state=s_tx_pdu_header;
						     r_crc_init=1'b1;
							 end
						
						  else
						    begin
							  r_tx_shift_reg=BLE_DATA_HEADER[15:0]; 
						     next_state=s_tx_pdu_header;
						     r_crc_init=1'b1;
							 end
												
						//状态机跳转时，把 r_crc_init 置为 1，即对 CRC 模块进行初始化；
		            //同时为了方便后续对数据载荷的提取，令 TX-RAM 的地址指针指向末尾处。		  
				   end
				 else next_state=s_tx_access; 
			  end
		   r_cnt=r_cnt+5'b1;		  
		  end
     s_tx_ci: //这个状态仅在发送报文为 1Mbps 编码类型时才会被用到 
	     begin
		    r_fsm_data=r_tx_shift_reg[0];
			 r_tx_shift_reg={1'b0, r_tx_shift_reg[31:1]};
			 if(r_cnt==5'd1) 
			   begin
					r_cnt=0;
					r_tx_shift_reg=BLE_TERM1[2:0]; 
				   next_state=s_tx_term1;
				end
			 else next_state=s_tx_ci;  
			 r_cnt=r_cnt+5'b1;	
		  end
     s_tx_term1: //这个状态在发送数据为 1Mbps 编码类型时才会被用到
	     begin
		    r_fsm_data=r_tx_shift_reg[0];
			 r_tx_shift_reg={1'b0, r_tx_shift_reg[31:1]};
			 if(r_cnt==5'd2)  //发送 3bits 的 TERM1，用来使 CODE 模块中的卷积编码器恢复初始状态
			   begin
					r_cnt=0;
					next_state=s_tx_pdu_header;
					if(BLE_ADV_STATE==0)  r_tx_shift_reg=BLE_ADV_HEADER[15:0]; 
					else                  r_tx_shift_reg=BLE_DATA_HEADER[15:0]; 
				end
			else next_state=s_tx_term1; 
			r_cnt=r_cnt+5'b1;
		  end
     s_tx_pdu_header: //公共部分
	     begin
		    r_fsm_data=r_tx_shift_reg[0];
			 r_tx_shift_reg={1'b0, r_tx_shift_reg[31:1]};
			 if(r_cnt==5'd1)  //r_cnt 计数到 1,把白化模块的使能信号置为有效状态，开始对 Header 部分进行白化操作。
			   begin
					r_switch_dwh=1;
					next_state=s_tx_pdu_header;
				end
			 else if(r_cnt==5'd11)
			   begin
		         RAM_A2=RAM_A2+7'b1;
					RAM_CS2=1;
					RAM_WEN2=0;
					RAM_OE2=1;
					PAYLOAD=0;
					next_state=s_tx_pdu_header;
			  //令 TX-RAM 的地址指针加 1，同时把 TX-RAM 的读使能信号置为有效状态，这样就可以从 TX-RAM中取出 32bits 的 payload
				end 
			 else if(r_cnt==5'd12)
			   begin
				   PAYLOAD=ram_d2;
					next_state=s_tx_pdu_header;
				end
			 else if(r_cnt==5'd15)
			   begin
					r_cnt=0;
					r_tx_shift_reg=PAYLOAD; 
				   next_state=s_tx_pdu_payload;
				end
			 r_cnt=r_cnt+5'b1;
		  end
     s_tx_pdu_payload: //公共部分
	     begin
		  //发送有效载荷部分，即 payload。
		    r_fsm_data=r_tx_shift_reg[0];
			 r_tx_shift_reg={1'b0, r_tx_shift_reg[31:1]};
		  //由于蓝牙设备可以发送不同长度的 payload，所以每次在 r_cnt 计数到 27 时，都会从 TX-RAM 中取出 32bits的 payload；
		    if(r_cnt==5'd7 && r_bytes==8'd1)
			  begin
               //RAM_CS2=0;
					RAM_OE2=0;
					next_state=s_wait_crc;
				 //从 TX-RAM 中取出 32bits的 payload
			  end
		    else if(r_cnt==5'd15 && r_bytes==8'd2)
			  begin
               //RAM_CS2=0;
					RAM_OE2=0;
					next_state=s_wait_crc;
				 //从 TX-RAM 中取出 32bits的 payload
			  end	
		    else if(r_cnt==5'd23 && r_bytes==8'd3)
			  begin
               //RAM_CS2=0;
					RAM_OE2=0;
					next_state=s_wait_crc;
				 //从 TX-RAM 中取出 32bits的 payload
			  end		  
			 else if(r_cnt==5'd27)
			  begin
			      RAM_A2=RAM_A2+7'b1;
               RAM_CS2=1;
					RAM_WEN2=0;
					RAM_OE2=1;
					next_state=s_tx_pdu_payload;
				 //从 TX-RAM 中取出 32bits的 payload
			  end
			 else if(r_cnt==5'd28)
			  begin
				   PAYLOAD=ram_d2;
					next_state=s_tx_pdu_header;
			  end
			 else if(r_cnt==5'd31)
			  begin
			      r_tx_shift_reg=PAYLOAD; 
					r_bytes=r_bytes-8'd4;
					r_cnt=0;
               if(r_bytes==0) 
					begin
					   r_cnt=0;
						next_state=s_wait_crc;
					end
					else next_state=s_tx_pdu_payload;
			  end
			 else next_state=s_tx_pdu_payload;
			 r_cnt=r_cnt+5'b1;
		  //在 r_cnt 计数到 31 时，把取出的 32bits payload 装入移位寄存器中，同时r_bytes 减 4。
		  //以此类推，直到 payload 全部发送完成，状态机才跳转至 s_wait_crc 状态，同时关闭该模块的输出使能信号。 
		  
		  //发送期间，用 r_bytes 指示 TX-RAM 中还有多少字节的 payload 没有被发送。
		  //如果设备发送报文中 payload 的长度为（4n+1）Bytes，则当 r_cnt 第（4n+1）次计数到7 时，发送完成。
		  //同理，payload 的长度为（4n+2）、（4n+3）、（4n+4）Bytes 时，当 r_cnt第（4n+1）次计数到 15, 23, 31 时，发送完成。 
        //next_state=s_wait_crc;
		  end
     s_wait_crc:  //公共部分
	     begin
		  //输出 24 个零给 CRC 模块，确保 24 位 CRC 码的发送。 
		   r_fsm_data=0;
         if(BLE_TYPE==3'b100) 
			  begin
			    if(r_cnt==5'd24)
				   begin
					   r_cnt=0;
						r_tx_shift_reg=BLE_TERM2[2:0];
						next_state=s_tx_term2;
				   end
				 else next_state=s_wait_crc;
				end
			else
			  begin
			    if(r_cnt==5'd24)
				   begin
					   r_cnt=0;
						next_state=s_end;
						tx_fsm_finished=1;
	     //状态机跳转到 s_end 状态时，表明状态机的发送已经完成，此时把 tx_fsm_finished置为有效状态并保持一个时钟周期，同时帧间隔计数器开始计数。
				   end
				 else next_state=s_wait_crc;
				end
		   r_cnt=r_cnt+5'b1;	
		  end
     s_tx_term2: 
	     begin
		  //当 TERM2 发送完成时，状态机跳转到 s_end 状态。这个状态仅在发送数据为 1M 编码类型时才会被用到。 
		    r_fsm_data=r_tx_shift_reg[0];
			 r_tx_shift_reg={1'b0, r_tx_shift_reg[31:1]};
			 if(r_cnt==5'd2)  //发送 3bits 的 TERM2，用来使 CODE 模块中的卷积编码器恢复初始状态。
			   begin
					r_cnt=0;
				   next_state=s_end;
				end
			 else next_state=s_tx_term2;
			 r_cnt=r_cnt+5'b1;
		  end
     s_end: 
	     begin
		  //此状态是为了给 PKA 模块中的的数据传送留出充足的时间，当把数据完整的发送出去之后，跳转到 s_reset 状态，同时把白化模块的使能信号置为无效状态。
		    next_state=s_reset;
			 r_switch_crc=0;
		  end		  
     s_reset: 
	     begin
		  //此状态是为了给 RIF 模块中的的数据传送留出充足的时间，当把数据完整的发送出去之后，跳转到 s_idle 状态。
		  //同时把 r_rst_tx 置为 1，用来关闭发送的时钟，并对一些信号进行初始化操作。 
          next_state=s_idle;
			 r_rst_tx_reg=1;
		  end	

	  default:
       begin
		   next_state=s_idle;
		 end
	  endcase
	  
	  //PAYLOAD=RAM_D;
 end
/*
 //当读使能有效，把所读数据读取到payload的寄存器中
 always@(RAM_REN)
  begin
   PAYLOAD=RAM_D;
  end
*/
 always@(posedge pka_1or2m_gck,negedge rst_n)
	if(!rst_n)
	 begin
	  current_state<=s_reset;
	 end
	else
	 current_state<=next_state;
	 //r_cnt<=r_cnt+5'b1;

endmodule